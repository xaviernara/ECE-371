library ieee;
use ieee.std_logic_1164.all;

entity btc_8bit is
  generic( SIGNED_OPS : boolean := true ); --(Un)signed feature
  port( x : in std_logic_vector(7 downto 0); --First operand
	y : in std_logic_vector(7 downto 0);  --Second operand
        z_GSE : out std_logic_vector(2 downto 0)--Comparison results 
	); 

end entity btc_8bit;

--The configurable BTC-8 operates on unsigned operands if feature parameter SIGNED_OPS = false
--and operates on signed two?s complement operands if feature parameter SIGNED_OPS = true. The
--BTC-8 comprises several CPC-2?s arranged in a binary tree. No other logic is allowed.
--
--In an architecture named structure, model the configurable BTC-8 using entity instantiation
--statements and named association. Also, use simple concurrent signal assignment statements and
--the concatenation operator. Additionally, consider using constant objects and the open keyword
--when appropriate.




architecture structure of btc_8bit is 

signal c1,c2,c3,c4,c5,c6,c7: std_logic_vector(2 downto 0);
constant un_signed : boolean := false;

begin

cpc_2bit1: entity work.cpc_2bit(dataflow)
 generic map(SIGNED_OPS=> SIGNED_OPS)
 port map(x=>x(7 downto 6),y=>y(7 downto 6),z_GSE=>c1);


cpc_2bit2: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map(x=>x(5 downto 4),y=>y(5 downto 4),z_GSE=>c2);
	

cpc_2bit3: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map(x=>x(3 downto 2),y=>y(3 downto 2),z_GSE=>c3);


cpc_2bit4: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map(x=>x(1 downto 0),y=>y(1 downto 0),z_GSE=>c4);
	
		
cpc_2bit5: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map(x=>c1(2) & c2(2),y=>c1(1) & c2(1),z_GSE=>c5);
	

cpc_2bit6: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map(x=>c3(2) & c4(2),y=>c3(1) & c4(1),z_GSE=>c6);
	

cpc_2bit7: entity work.cpc_2bit(dataflow)
generic map(SIGNED_OPS=> un_signed)
port map (x=>c5(2) & c6(2),y=>c5(1) & c6(1),z_GSE=>c7);

z_GSE<=c7;

end architecture structure;
		