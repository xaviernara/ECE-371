library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity p3_fetch_no_bypass is
	generic (SIZE : positive :=32);
	port(Branch_Mux_Control_RT_GSED: in std_logic_vector(1 downto 0); --FROM CONTROL UNIT
		WREN,clk,rst : IN std_logic;
		BTA_IN_FETCH : IN std_logic_vector(31 downto 0);
		JRTA_IN_FETCH : IN std_logic_vector(31 downto 0);
		JTA_IN_FETCH : IN std_logic_vector(31 downto 0);
		DATA : in std_logic_vector(31 downto 0);
		CLA_COUT_PC_PLUS_1 : OUT std_logic;
		CLA_Y_PC_PLUS_1 : in std_logic_VECTOR (7 DOWNTO 0);
		CLA_sum_out : OUT std_logic_vector(7 downto 0);


		rd1inein_DECODE : out std_logic_vector(31 downto 0);
		PC1in_DECODE : out std_logic_vector(31 downto 0)
	);
end entity p3_fetch_no_bypass;

architecture structure of p3_fetch_no_bypass is

	signal ADD_INSTRUCTION: std_logic_vector(31 downto 0);
	signal rd1ineout_FETCH : std_logic_vector(31 downto 0);
	signal PC1out_FETCH : std_logic_vector(31 downto 0);
	signal INSTRUCTION_ADD_OUT : std_logic_vector(31 downto 0);
	signal PC_Plus1 : std_logic_vector(31 downto 0);
	--signal CLA_sum_out : std_logic_vector(7 downto 0);
	--signal PCPLUS_1_cout : std_logic_vector(7 downto 0);

begin

--PC + 1 SECTION
PC_PLUS1<= INSTRUCTION_ADD_OUT or 32x"1";
PC1out_FETCH <= PC_Plus1;

Instruction_Memory : entity work.instructionROM(SYN)
	generic map(SIZE => SIZE )
	port map(aclr => '0', address => ADD_INSTRUCTION(7 downto 0) ,clken => '1' ,clock => clk, data=>DATA, wren=>WREN, q => rd1ineout_FETCH );


SELECT_Address: entity work. mux_4to1(behavhior)
	generic map (SIZE=> SIZE)
	port map (w0 => PC_Plus1, w1 => JRTA_IN_FETCH, w2 => BTA_IN_FETCH, w3 => JTA_IN_FETCH, s => Branch_Mux_Control_RT_GSED, f => ADD_INSTRUCTION);

CLA_PC_PLUS_1: ENTITY work. cla_8bit(structure)
port map (x=>PC1out_FETCH(31 DOWNTO 24) ,y=>CLA_Y_PC_PLUS_1,cin=>'0',cout=>CLA_COUT_PC_PLUS_1 ,sum=>PC_PLUS1(31 DOWNTO 24),GG =>OPEN,GA =>OPEN);



----------------------------------------------------------------------------------------------------------------------------
------------------------------------------------------Through the pipeline (ie the output signals going thru to the decode STAGE)--------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------

	d_FLIP_flopforPC1 : entity work.dflop(behavior)
			generic map(SIZE=>SIZE)
			port map(clk => clk, rst => rst, clken => '1', din => PC1out_FETCH, q => PC1in_DECODE);

	d_FLIP_flopforRD : entity work.dflop(behavior)
			generic map(SIZE=>SIZE)
			port map(clk => clk, rst => rst, clken => '1', din => rd1ineout_FETCH, q => rd1inein_DECODE);

	d_FLIP_flopBEFOREPC1: entity work.dflop(behavior)
			generic map(SIZE=>SIZE)
			port map(clk => clk, rst => rst, clken => '1', din =>  ADD_INSTRUCTION, q => INSTRUCTION_ADD_OUT );


END ARCHITECTURE STRUCTURE;

	